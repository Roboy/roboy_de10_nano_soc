// soc_system_auxilliary.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module soc_system_auxilliary (
		input  wire [3:0]  I2C_0_avalon_slave_0_address,     // I2C_0_avalon_slave_0.address
		input  wire        I2C_0_avalon_slave_0_write,       //                     .write
		input  wire [31:0] I2C_0_avalon_slave_0_writedata,   //                     .writedata
		input  wire        I2C_0_avalon_slave_0_read,        //                     .read
		output wire [31:0] I2C_0_avalon_slave_0_readdata,    //                     .readdata
		output wire        I2C_0_avalon_slave_0_waitrequest, //                     .waitrequest
		input  wire        I2C_0_clock_sink_clk,             //     I2C_0_clock_sink.clk
		inout  wire        I2C_0_conduit_end_scl,            //    I2C_0_conduit_end.scl
		inout  wire        I2C_0_conduit_end_sda,            //                     .sda
		input  wire        I2C_0_reset_reset,                //          I2C_0_reset.reset
		input  wire [3:0]  I2C_1_avalon_slave_0_address,     // I2C_1_avalon_slave_0.address
		input  wire        I2C_1_avalon_slave_0_write,       //                     .write
		input  wire [31:0] I2C_1_avalon_slave_0_writedata,   //                     .writedata
		input  wire        I2C_1_avalon_slave_0_read,        //                     .read
		output wire [31:0] I2C_1_avalon_slave_0_readdata,    //                     .readdata
		output wire        I2C_1_avalon_slave_0_waitrequest, //                     .waitrequest
		input  wire        I2C_1_clock_sink_clk,             //     I2C_1_clock_sink.clk
		inout  wire        I2C_1_conduit_end_scl,            //    I2C_1_conduit_end.scl
		inout  wire        I2C_1_conduit_end_sda,            //                     .sda
		input  wire        I2C_1_reset_reset,                //          I2C_1_reset.reset
		input  wire [3:0]  I2C_2_avalon_slave_0_address,     // I2C_2_avalon_slave_0.address
		input  wire        I2C_2_avalon_slave_0_write,       //                     .write
		input  wire [31:0] I2C_2_avalon_slave_0_writedata,   //                     .writedata
		input  wire        I2C_2_avalon_slave_0_read,        //                     .read
		output wire [31:0] I2C_2_avalon_slave_0_readdata,    //                     .readdata
		output wire        I2C_2_avalon_slave_0_waitrequest, //                     .waitrequest
		input  wire        I2C_2_clock_sink_clk,             //     I2C_2_clock_sink.clk
		inout  wire        I2C_2_conduit_end_scl,            //    I2C_2_conduit_end.scl
		inout  wire        I2C_2_conduit_end_sda,            //                     .sda
		input  wire        I2C_2_reset_reset,                //          I2C_2_reset.reset
		input  wire [3:0]  I2C_3_avalon_slave_0_address,     // I2C_3_avalon_slave_0.address
		input  wire        I2C_3_avalon_slave_0_write,       //                     .write
		input  wire [31:0] I2C_3_avalon_slave_0_writedata,   //                     .writedata
		input  wire        I2C_3_avalon_slave_0_read,        //                     .read
		output wire [31:0] I2C_3_avalon_slave_0_readdata,    //                     .readdata
		output wire        I2C_3_avalon_slave_0_waitrequest, //                     .waitrequest
		input  wire        I2C_3_clock_sink_clk,             //     I2C_3_clock_sink.clk
		inout  wire        I2C_3_conduit_end_scl,            //    I2C_3_conduit_end.scl
		inout  wire        I2C_3_conduit_end_sda,            //                     .sda
		input  wire        I2C_3_reset_reset                 //          I2C_3_reset.reset
	);

	I2C_avalon_bridge #(
		.CLOCK_SPEED_HZ (50000000),
		.BUS_SPEED_HZ   (400000)
	) i2c_0 (
		.reset       (I2C_0_reset_reset),                //          reset.reset
		.address     (I2C_0_avalon_slave_0_address),     // avalon_slave_0.address
		.write       (I2C_0_avalon_slave_0_write),       //               .write
		.writedata   (I2C_0_avalon_slave_0_writedata),   //               .writedata
		.read        (I2C_0_avalon_slave_0_read),        //               .read
		.readdata    (I2C_0_avalon_slave_0_readdata),    //               .readdata
		.waitrequest (I2C_0_avalon_slave_0_waitrequest), //               .waitrequest
		.scl         (I2C_0_conduit_end_scl),            //    conduit_end.scl
		.sda         (I2C_0_conduit_end_sda),            //               .sda
		.clock       (I2C_0_clock_sink_clk)              //     clock_sink.clk
	);

	I2C_avalon_bridge #(
		.CLOCK_SPEED_HZ (50000000),
		.BUS_SPEED_HZ   (400000)
	) i2c_1 (
		.reset       (I2C_1_reset_reset),                //          reset.reset
		.address     (I2C_1_avalon_slave_0_address),     // avalon_slave_0.address
		.write       (I2C_1_avalon_slave_0_write),       //               .write
		.writedata   (I2C_1_avalon_slave_0_writedata),   //               .writedata
		.read        (I2C_1_avalon_slave_0_read),        //               .read
		.readdata    (I2C_1_avalon_slave_0_readdata),    //               .readdata
		.waitrequest (I2C_1_avalon_slave_0_waitrequest), //               .waitrequest
		.scl         (I2C_1_conduit_end_scl),            //    conduit_end.scl
		.sda         (I2C_1_conduit_end_sda),            //               .sda
		.clock       (I2C_1_clock_sink_clk)              //     clock_sink.clk
	);

	I2C_avalon_bridge #(
		.CLOCK_SPEED_HZ (50000000),
		.BUS_SPEED_HZ   (400000)
	) i2c_2 (
		.reset       (I2C_2_reset_reset),                //          reset.reset
		.address     (I2C_2_avalon_slave_0_address),     // avalon_slave_0.address
		.write       (I2C_2_avalon_slave_0_write),       //               .write
		.writedata   (I2C_2_avalon_slave_0_writedata),   //               .writedata
		.read        (I2C_2_avalon_slave_0_read),        //               .read
		.readdata    (I2C_2_avalon_slave_0_readdata),    //               .readdata
		.waitrequest (I2C_2_avalon_slave_0_waitrequest), //               .waitrequest
		.scl         (I2C_2_conduit_end_scl),            //    conduit_end.scl
		.sda         (I2C_2_conduit_end_sda),            //               .sda
		.clock       (I2C_2_clock_sink_clk)              //     clock_sink.clk
	);

	I2C_avalon_bridge #(
		.CLOCK_SPEED_HZ (50000000),
		.BUS_SPEED_HZ   (400000)
	) i2c_3 (
		.reset       (I2C_3_reset_reset),                //          reset.reset
		.address     (I2C_3_avalon_slave_0_address),     // avalon_slave_0.address
		.write       (I2C_3_avalon_slave_0_write),       //               .write
		.writedata   (I2C_3_avalon_slave_0_writedata),   //               .writedata
		.read        (I2C_3_avalon_slave_0_read),        //               .read
		.readdata    (I2C_3_avalon_slave_0_readdata),    //               .readdata
		.waitrequest (I2C_3_avalon_slave_0_waitrequest), //               .waitrequest
		.scl         (I2C_3_conduit_end_scl),            //    conduit_end.scl
		.sda         (I2C_3_conduit_end_sda),            //               .sda
		.clock       (I2C_3_clock_sink_clk)              //     clock_sink.clk
	);

endmodule
